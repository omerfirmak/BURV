module lsu (
	input clk,    // Clock
	input rst_n   // Asynchronous reset active low
	
);

endmodule